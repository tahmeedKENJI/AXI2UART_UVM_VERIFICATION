`ifndef _DEPENDENCIES_SVH_
`define _DEPENDENCIES_SVH_

`include "uvm_macros.svh"
import uvm_pkg::*;

`endif

